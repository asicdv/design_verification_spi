/*
 * Author:  Deepak Siddharth Parthipan
 *          RIT, NY, USA
 * Module:  Package
 */
//-------------------------------------------------------------
package spi_pkg;
//-------------------------------------------------------------
	import uvm_pkg::*;

    //`include "uvm_macros.svh"
    `include "spi_tb_defines.sv"
    `include "spi_sequence_item.sv"
	`include "spi_driver.sv"
	`include "spi_monitor.sv"
	`include "spi_sequencer.sv"
	`include "spi_agent.sv"
	`include "spi_scoreboard.sv"
    `include "spi_sequence.sv"
	`include "spi_env.sv"
	`include "spi_test.sv"
//-------------------------------------------------------------
endpackage: spi_pkg
//-------------------------------------------------------------
